module DE10_lite_switch_controller(
    input clk,

    input [9:0] sw_toggle,
    input [9:0] sw_out
);





endmodule